���Z     @  L   I     �  &                                       
    �                                                    !   �   �V 	   ,          � Project@Options� -�   !�     7   \+ 	   -          � File@@Version2.1  � 1.1     (                                                          1   f   TOPIC VERSION OBJARRAY BROWSE_SEQUENCE BUILD_TAG CONTEX    link viewHandles 7                                            _ISECT_iterator _AE_Sorter _AE_mark _SysInfoFlags _outside_   Metafile VbPicture VbVarArray VeRec ViewEngine WinImage _AE   r VB_Historian VB_View VbCurrency VbDibBitmap VbFixArray Vb	   ng SystemDatabase TextFileDatabase TrashCollector TreeWalke
   Real RecordMark RuleSpecifier SchemaEngine SmartString Stri   adStream NamedData NamedMonad NilMonad Number Presentation    Dictionary Integer LogStream Monad MonadArray MonadFile Mon   tion Bcd36 Boolean ClassDesc ClassMethod ComboElement Date    Set AdRec AeAccessSet AgilityDatabase ArrayDatabase Associa   ]  YAccessCombo AccessEngine AccessItem AccessRule Access`, �                  .       ,       )       Q       �     :�     �L     ��     ��     ��     ��     ��     ��     �4     ��     �!     �/     �)     �     �     ��     ��     �L     `     M     `     Fx     r     ��     ��     ��     ��     ��     �     ��     ��     ��     ��     �1     �<     ��     �?      ��     ��     ��     �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �0    !� BuildAll!� 0!� Contents!� Copyright � pi & alex!�  #     �  �� 	\�   O -�   !� /T N /Just L /Text ������!� /Z     N /Style /Just L!� /X /Style /Just L  
q �              F   ,192), 0!�3 "Index", ( 511, 0, 511, 1023), , , (192,192,192$   192,192), 0!�4 "Glossary", ( 0, 0, 511, 1023), , , (192,192%   , , (192,192,192), 0!�. "", ( 0, 511, 1023, 511), , , (192,&   832, 832), , , (192,192,192), 0!�, "", ( 0, 0, 1023, 511), '   ' "Visual Expert", , , , (192,192,192), 0!�- "", ( 64, 64, (   �  �� 	   -          � F1ProjectWindowso-�  � !�    �  !�  !�  !�  !�  !�                                      *     !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !+   �   �� 	   -          � F1ProjectButtonsZ -�   !��  �, "����� �����",(Global), 0,<Dlg_FolderSelect>!� ��������-   0  � 	   .          � F1ProjectGlossary -�  # !    No!�  !� Visual Expert!� 1!�  !�  !�  !�                 /   !�  !� F:\WORK\expert\rc\vs.ico!� 0!�  !�  !� 0!� 0!� �    T_STRING HELP_MACRO KEYWORDS TOPIC_TITLE NOTE              >   ay /popup/Text ������L�L, /Jump Window_All /Link /Macro /P4   ������� - ��������� ������ �������� ������ � ������� ��. ��5   �� �� ����, �� ��������� ����� �������. ����� ��������� ���   �� ���������� ��.!�2 /S /Just L /Text ������ �����  ������ 1  ������������� V�     �  �� 	fM  �-�   !�  /T N /JustO  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !� 9  ork\expert\hlp\close.bmp /Macro /Play /Popup /Just L  
� 8   ext ������ ����� ������ ������������!�G /I /Jump /Link f:\wE   �� ��L�L, /Jump Window_All /Link /Macro /Play /popup/Text:   �L�L, /Jump Window_All /Link /Macro /Play /popup/Text �����;   /Jump Window_All /Link /Macro /Play /popup/Text �����������<   l /Link /Macro /Play /popup/Text ������� �������������L�L, =   lay /popup/Text ������� ���������������L�L, /Jump Window_Al@   �   �'�� 
� ( / D     � Topic@Index  �    �  "     �    �  ��6S     �  �� =h   
  � Index�� Lx   6H   � ������L�L, /Jump Admin_Admin /Link /Macro /Play /popup/T@  ���� �������L�L, /Jump HelpHlp /Link /Macro /Play /popup/TB   t �������L�L, /Jump HelpHlp /Link /Macro /Play /popup/Text C   opup/Text ���������� ����B�B,/Link /Macro /Play /Popup/TexD    ��������� ����L�L, /Jump Window_All /Link /Macro /Play /pJ   ), 0!�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !� 2   �� ���������� ������L�L, /Jump Window_All /Link /Macro /PlG   ext �����������������B�B,/Link /Macro /Play /Popup/Text ��  ���� ������������!�^ /L /Jump Protect /Link /Macro /Play /p%   !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  ���� � ��������� �������� Visual Expert�!�1 /S /Just L /TexM   �������� ������������ � ������� ���� ���������� ���������� N   ������.!�� /B /Just L /Text ����� �������������� �� � ����O   ��� �������� ������ ��� �����. ��� ������ ������ ������ ���K   ���� ��� ��� �������� ���������� ��, ������� ������ ������    , !�                                                       `   0'  y. 	   ,          � F1ProjectStyle2'-�  � !�Ha   0 , None , !�H Heading , Arial ,  12 ,  180 ,  250 ,  60 , R   ding , System ,  12 ,  180 ,  250 ,  60 ,  20 ,  0 , -1 ,  S   0 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�I HeaT   20 ,  60 ,  0 ,  0 ,  0 , None , !�J Paragraph , Arial ,  1U   ,  0 , None , !�J Paragraph , Arial ,  10 ,  180 ,  250 ,  V   aragraph , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 W    10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�J PX     20 ,  60 ,  0 ,  0 ,  0 , None , !�J Paragraph , Arial , Y    ,  0 , None , !�K Paragraph , System ,  10 ,  180 ,  250 ,Z   !�F Title , Arial ,  18 ,  120 ,  250 ,  40 ,  40 ,  0 , -1[   al ,  18 ,  120 ,  250 ,  40 ,  40 ,  0 , -1 ,  0 , None , \    ,  250 ,  40 ,  40 ,  0 , -1 ,  0 , None , !�F Title , Ari]     40 ,  0 , -1 ,  0 , None , !�F Title , Arial ,  18 ,  120^     0 , Shade , !�F Title , Arial ,  18 ,  120 ,  250 ,  40 ,_    Title , System ,  18 ,  120 ,  250 ,  40 ,  40 ,  1 , -1 ,�p    20 ,  0 , -1 ,  0 , None , !�H Heading , Arial ,  12 ,  18q     0 , None , !�L Jump Label , Arial ,  10 ,  180 ,  250 ,  b    Label , Arial ,  10 ,  180 ,  250 ,  20 ,  20 ,  10 ,  0 ,c   ,  180 ,  250 ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�L Jumpd     20 ,  10 ,  0 ,  0 , None , !�L Jump Label , Arial ,  10 e    None , !�M Jump Label , System ,  10 ,  180 ,  250 ,  20 ,f   ng , Arial ,  12 ,  180 ,  250 ,  40 ,  20 ,  0 , -1 , -1 ,g   80 ,  250 ,  40 ,  20 ,  0 , -1 , -1 , None , !�L Sub Headih    ,  0 , -1 , -1 , None , !�L Sub Heading , Arial ,  12 ,  1i   e , !�L Sub Heading , Arial ,  12 ,  180 ,  250 ,  40 ,  20j    Arial ,  12 ,  180 ,  250 ,  40 ,  20 ,  0 , -1 , -1 , Nonk     250 ,  40 ,  20 ,  1 , -1 , -1 , None , !�L Sub Heading ,l    , -1 ,  0 , None , !�M Sub Heading , System ,  12 ,  180 ,m    , !�H Heading , Arial ,  12 ,  180 ,  250 ,  60 ,  20 ,  0n   Arial ,  12 ,  180 ,  250 ,  60 ,  20 ,  0 , -1 ,  0 , Noneo   0 ,  250 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�H Heading ,    20 ,  20 ,  10 ,  0 ,  0 , None , !�L Jump Label , Arial , �   ,  0 ,  0 , None , !�S Bitmap Paragraph , System ,  18 ,  1r   , !�H Footnote , Arial ,  8 ,  180 ,  250 ,  20 ,  60 ,  0 s   Arial ,  8 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None t    ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�H Footnote , u   60 ,  0 ,  0 ,  0 , None , !�H Footnote , Arial ,  8 ,  180v    , None , !�H Footnote , Arial ,  8 ,  180 ,  250 ,  20 ,  w   note , System ,  8 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0x    ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�I Footy    60 ,  0 ,  0 ,  0 , None , !�N Mono Spaced , Courier ,  10z   ne , !�N Mono Spaced , Courier ,  10 ,  180 ,  250 ,  20 , {   Courier ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , No|    250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�N Mono Spaced , }     0 ,  0 , None , !�N Mono Spaced , Courier ,  10 ,  180 , ~   Mono Spaced , System ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,    10 ,  180 ,  250 ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�M    80 ,  250 ,  20 ,  60 ,  1 , -1 ,  0 , Shade , !�Q Bitmap P�    , None , !�G Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  6�   let , System ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0�   0 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�H Bul�    ,  0 ,  0 ,  0 , None , !�R Bitmap Jump Label , Arial ,  1�   R Bitmap Jump Label , Arial ,  10 ,  180 ,  250 ,  20 ,  60�    ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !��   ,  60 ,  0 ,  0 ,  0 , None , !�R Bitmap Jump Label , Arial�    , !�R Bitmap Jump Label , Arial ,  10 ,  180 ,  250 ,  20 �   stem ,  10 ,  180 ,  250 ,  20 ,  60 ,  10 ,  0 ,  0 , None�   20 ,  60 ,  0 ,  0 ,  0 , None , !�T Bitmap Jump Label , Sy�   None , !�Q Bitmap Paragraph , Arial ,  10 ,  180 ,  250 ,  �   h , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , �   250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�Q Bitmap Paragrap�   ,  0 , None , !�Q Bitmap Paragraph , Arial ,  10 ,  180 ,  �   aragraph , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0     0 ,  0 ,  0 ,  0 , None , !�G Bullet , Arial ,  10 ,  180 ,�    250 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�M Outline Node ,�   ,  0 ,  0 , None , !�M Outline Node , Arial ,  10 ,  180 , �    Outline Node , Arial ,  10 ,  180 ,  250 ,  10 ,  10 ,  0 �   ,  10 ,  180 ,  250 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�M�   20 ,  60 ,  0 ,  0 ,  0 , None , !�N Outline Node , System �   one , !�R Enumerated Bullet , Arial ,  10 ,  180 ,  250 ,  �    , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , N�   0 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�R Enumerated Bullet�   0 , None , !�R Enumerated Bullet , Arial ,  10 ,  180 ,  25�   ullet , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  �   ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�R Enumerated B�    ,  0 , None , !�S Enumerated Bullet , System ,  10 ,  180 �   �G Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0�   l ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�     250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�G Bullet , Aria��    Arial ,  10 ,  180 ,  250 ,  10 ,  10 ,  0 ,  0 ,  0 , Non�    ,  60 ,  0 ,  0 ,  0 , None , !�T Index Letter Label , Sys�    0 ,  0 , None , !�E Line , Arial ,  10 ,  180 ,  250 ,  20�    , !�E Line , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 , �   Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None�    180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�E Line , �    20 ,  60 ,  0 ,  0 ,  0 , None , !�E Line , Arial ,  10 , �   ,  0 ,  0 , None , !�F Line , System ,  10 ,  180 ,  250 , �    Outline Leaf , Arial ,  10 ,  440 ,  250 ,  10 ,  10 ,  0 �   ,  10 ,  440 ,  250 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�M�    10 ,  10 ,  0 ,  0 ,  0 , None , !�M Outline Leaf , Arial �    0 , None , !�M Outline Leaf , Arial ,  10 ,  440 ,  250 , �   e Leaf , Arial ,  10 ,  440 ,  250 ,  10 ,  10 ,  0 ,  0 , �     440 ,  250 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�M Outlin�   0 ,  0 ,  0 ,  0 , None , !�N Outline Leaf , System ,  10 ,�   e , !�M Outline Node , Arial ,  10 ,  180 ,  250 ,  10 ,  16�   tem ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , None ,�   tter Label , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -�    ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , None , !�V Glossary Le�    0 , None , !�W Glossary Letter Label , System ,  12 ,  180�    Index , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 , �   ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F�    250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Index , Arial �   0 ,  0 ,  0 ,  0 , None , !�F Index , Arial ,  10 ,  180 , �   0 , None , !�F Index , Arial ,  10 ,  180 ,  250 ,  20 ,  6�   ndex , System ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  �    12 ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , None , !�G I�   0 ,  0 , -1 ,  0 , None , !�S Index Letter Label , Arial , �   S Index Letter Label , Arial ,  12 ,  180 ,  250 ,  20 ,  6�    ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , None , !��     60 ,  0 , -1 ,  0 , None , !�S Index Letter Label , Arial�    !�S Index Letter Label , Arial ,  12 ,  180 ,  250 ,  20 ,��   1 ,  0 , None , !�V Glossary Letter Label , Arial ,  12 ,  �    , None , !�F Image , Arial ,  10 ,  180 ,  250 ,  20 ,  60�   mage , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0�    10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F I�   50 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Image , Arial , �     0 ,  0 ,  0 , None , !�G Image , System ,  10 ,  180 ,  2�   ne , !�I Glossary , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,�   , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , No�   80 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�I Glossary �    60 ,  0 ,  0 ,  0 , None , !�I Glossary , Arial ,  10 ,  1�    , None , !�I Glossary , Arial ,  10 ,  180 ,  250 ,  20 , �   ary , System ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0�   ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , None , !�J Gloss�   , -1 ,  0 , None , !�V Glossary Letter Label , Arial ,  12 �    Letter Label , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 �   180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , None , !�V Glossary�    ,  0 ,  0 ,  0 , None , !�F Image , Arial ,  10 ,  180 ,  �    None , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  �   e , !�;  , Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,�    Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , Non�    180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Table ,�   20 ,  60 ,  0 ,  0 ,  0 , None , !�F Table , Arial ,  10 , �     0 ,  0 , None , !�F Table , Arial ,  10 ,  180 ,  250 ,  �    , !�F Table , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,�   ystem ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None�   80 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�G Table , S�   20 ,  60 ,  0 ,  0 ,  0 , None , !�D Bar , Arial ,  10 ,  1�    ,  0 ,  0 , None , !�D Bar , Arial ,  10 ,  180 ,  250 ,  �   None , !�D Bar , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0�   r , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , �   10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�D Ba�   250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�D Bar , Arial ,  b�   , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1 �   ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  �    !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  �   None , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  ,�    , !�;  , Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , �     0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , �   ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,�    ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 �    0 ,  0 ,  0 ,  0 , None , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0�    0 ,  0 ,  0 ,  0 ,  , !�;  , Arial ,  10 ,  0 ,  0 ,  0 , �     0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 , �   ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,�    ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 �   10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�1  ,  ,  0�    0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�;  , Arial ,  �    ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,    0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�;  , Arial ,  1   ������������� ������ (�������� ����), � ���������� ������   ������������!�F /I /Jump /Link f:\work\expert\hlp\open.bmp I   rface /Link /Macro /Play /popup /Just L /Text ������ �������   rt\rc\yes.bmp /Just M /Text ����������!�] /L /Jump UserInte�   � P�     �  �� 	`}  �-�   !�= /R N /Link f:\work\expe�      � 0   �  ��9W     �  �� Aq     �
 �����������P    0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  �     0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , �   ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,�   0 ,  0 ,  0 ,  0 , None , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 �   0 ,  0 ,  0 ,  0 ,  , !�;  , Arial ,  10 ,  0 ,  0 ,  0 ,  �    0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  �     0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 , �   ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,�   0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�1  ,  ,  0 �  �� (������� ������ �����������).!�1 /S /Just L /Text ������  opup /Just L /Text ������ ������ � ������������� �������!�J  ��!�# /B /Just L /Text ������������� ����!�+ /S /Just L /Te  xt ������ �� ���������������:!� /B /Just L /Text ����� ���  ���.!�1 /B /Just L /Text ������ ����� � ������� ��������.      
 �                                                     ?  ���!�� /P /Just L /Text ��������� �������� ����� ���� �����  -�   !�4 /T N /Just M /Text ��������� �������� ������ ����  ������� �������� ������ ��������� Z�     �  �� 	j�  		     �  	  � 3020   �  ��@a     �  �� K�   &  �! ��  �  ���� 
� , 3 L     � Topic@File_Exit  �    �    	  � 3007   �  ��:[     �  �� Ez     � ����� ��   �������� T�     �  �� 	d�  ?-�   !� /T N /Just M /�  Text �����!�� /P /Just L /Text ���������� ����������. ��� �    \hlp\save.bmp /Macro /Play /Popup /Just L  
� �             ����� ������ ������������!�F /I /Jump /Link f:\work\expert�    /L /Jump MenuCommands /Link /Macro /Play /popup /Just L /T   ��������L�L, /Jump File_Recent /Link /Macro /Play /popup/T  ext ��������� �������� ������L�L, /Jump File_Exit /Link /Ma  cro /Play /popup/Text �����B�B,/Link /Macro /Play /Popup/T  ext �����������������L�L, /Jump Admin_ChangeLvl /Link /Mac  ro /Play /popup/Text �������� ������� ��������L�L, /Jump AdA   min_ChangeLvl /Link /Macro /Play /popup/Text ������� ������    /Macro /Play /Popup /Just L  
� �                        ^  ��� � ������������� ��������� R�     �  �� 	bk  �-�  Z  ��� ������� �� ������:  ������������, ����������� ���������z  ����� ������� ���������� (� �������� ������) ��� ����������H  ��!�M /K /Jump /Link /Macro /Play /Popup /Just L /Text ����_  lay /popup /Just L /Text ���������� �� �������� �����������  �, ������������� ������!�k /L /Jump FuncToc /Link /Macro /P  /Just L /Text ������������� ������, ���������� ������ �����  ext ������� ����!�y /L /Jump LL1 /Link /Macro /Play /popup   ��������L�L, /Jump File_Save /Link /Macro /Play /popup/Text#  ����� ��������� ������ ������ � ������������� �������. ����>  ������ ������, ���������� ��� �������� ��� ������� � ������7   �  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  $    !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !    ����� ����� ������ ������� ��.  
� �                     &  �������� � ������ ��������� �������������� ��. ����� ���� �'  L /Text ��� �������� ���� �� ����� �� ������-������������ �(  �+ /T N /Just M /Text ��������� �������� �����!�� /P /Just )  ��� �������������� ������� V�     �  �� 	f|  � -�   !,  �� ������ W�     �  �� 	g�  �-�   !� /T N /Just M /-  Text ������� ����!��/O /Just L /Cols 1 /Rows 22 /Type O /T.  ext B�B,/Link /Macro /Play /Popup/Text ����L�L, /Jump File/  _NewES /Link /Macro /Play /popup/Text ����� ���������� ����0  ����L�L, /Jump File_Open /Link /Macro /Play /popup/Text ���!  �����L�L, /Jump File_Save /Link /Macro /Play /popup/Text ��b"   M /Text �������������!�� /P /Just L /Text ��������� ������A  ����� ����� ������ ������������!�H /I /Jump /Link f:\work\e2  ��� ������������ �� ������� ��������.!�1 /S /Just L /Text �5    ���� 
� * 1 F     � Topic@HotKeys  �    �  6    �    �  ��8U     �  �� ?l     � HotKeys�� N|7       �  �� 	^   -�   !�+ /T N /Just M /Text ������� �(  ������� �������!�F /I /Jump /Link f:\work\expert\hlp\keys.w6    �  	  � 3022   �  ��<]     �  �� G~     � ������    �                                                          ;  ��� ��������� ������. � ������ ������ �������� ���� � ���� 9   ��� ������� ������ ��������� ������������.!�1 /S /Just L /T�   �  �a�� 
� + 2 H     � Topic@Contents  �    � �    � ������ ��������� (�� ��������� ��), �� ����� ������� ���  ��� ��������:!�C /K /Jump Dlg_Adm_Acc /Link /Macro /Play /p�  ������������. ��������_�������_������� ��� ������ ���������    ext ��������� �������  
� �                              �P  xpert\hlp\window.bmp /Macro /Play /Popup /Just L!�| /P /JusC  ��������� U�     �  �� 	e�  $-�   !�! /T N /Just M /'  Text ������ �������!�` /P /Just L /Text ������� ��������� ��  ��� �����. ����� �� ������ ����� �� ������� Esc.!�G /I /JumD  � ���� ����� ������� ���� ���������� ������� � ������������E  ���� ����� ������� � ��������� �������� ����. ����� �������F  ��� ��������� ������. � ���� ������ ������ ���� ��������� �K  ���� ������������� �����!�g /K /Jump Work /Link /Macro /Pla�   ���� ����� ����.!�s /K /Jump Admin_ChangeLvl /Link /Macro   �� ��� ������!�'/P /Just L /Text �������� MDI-���� ����� �J  y /popup /Just L /Text ������ ��������/�������� �����������M  �  [u�� 
� / 6 O     � Topic@MenuCommands  �  +    �  	  � 3000   �  ��=^     �  �� Hz     � ������  �������� ���� ����������� ������������� �� ��������� ����.�   !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�N  t L /Text ����� ������ ������������ �������� ���� - ������ �B  �  	  � 3050   �  ��;\     �  �� Fz     � ������ a  ���� ������ ���������, �� �������� ������ �����������.�����R  ����. ��������, ������� ������������ �������� �� ����� ����S  �� ������� ������������ ��� ������ ������������� ���� �� ��T   ����������. ���������� ������������ ������ ������������� �U   ��������� ������ � �������� ������� � ����� ������ �������V  ���������� ������������� ����-��� ������ ����. ������ �����W  ����� ����������. ������ ������������ ����� ������. ��� ���X  ����������, �������������. ��� ����������� � ������� ������Y  ���, �������, ����������� �������, ����������, �����������   y /Popup /Just L!��/P /Just L /Text ���  ������������ ����[  ��!�E /I /Jump /Link f:\work\expert\hlp\acc.wmf /Macro /Pla\  ���!�6 /H /Just L /Text ������������� ������� � ������ ����]   !�8 /T N /Just M /Text ������ ������ � ������������� ����I  ������ �� ��������� ������� - ������ ����� ������ ���������Q  �  ́�� 
 - 4 M     � Topic@StatusLine  �    bp   �������� ����������� ������� ��� ������������� ������� ���c  ����������������� � ������������ ��� �������� �� ��������, d  �������������� � ������������� ���������� ������ � ��������e  � ������. ���� ����� ���������� � ����� �� ���������� �����f  ���� ������ �� ������� ������������� ��� ������ (����������g  ���� ��� �������������) ����� �� ��������� �������. �������h  ��� ��������� �������������:!�U /K /Jump Explorer /Link /Mai  cro /Play /popup /Just L /Text ��������� ���������� ������!j  �u /K /Jump ProductEdit /Link /Macro /Play /popup /Just L /  Text �������� ������������� ��� ������, ��� �������� � ����    ���� - ������������� ������������.  
� �                 k  ��� ����� � ����� ��������������� ����������� ������ ������l  ������� � ������ ������� ����������.��!�n /P /Just L /Text m  �������� �������������. �� � ������ ������ ��������� ������n  �� ����� �������� � ������ ������� ����� ������� ������ ���o  ���� ���������� (�������� ������). � ���������� �����������b  � ��������� ������ ����������� � ���� ����. �������� ���� ��  e /Link /Macro /Play /popup /Just L /Text ������ �������!�Jr  ����� ������������ �������� MDI-����.!�J /K /Jump StatusLins  ������ ������� ���������� ������ �������� ����� ��������� �t  �������� ��������� ������ � ���. �������� �������� ��� ����u  , �� ��� ��������, ��������� ����� ������� ���� ������ ����v  �� ��������������/������������� �������� ���������� �������w  ������ �������� ������ ����������. ��������� ������� ������x  ������� ������ ��� �������� ������� � �������� ����� ������y   ����� �������. ���������� ������ ������������ ���������� �|  ����� �������������� X�     �  �� 	h�  -�  	 !�4 /T }  N /Just M /Text ��������� ���������� ������������!�p/P /Ju~  st L /Text ���������� ����� ���������������� ��������� ����  ����� �� ������������� ������ ���� - "���� ���������� ������  ��". ������ �������� ���� ������������� ����� ���������� ��q  ����� � ��� ��������� �������������� � ������������� �� � ��   /K /Jump MenuCommands /Link /Macro /Play /popup /Just L /T�   M /Text ��������� ����� � �����!�� /P /Just L /Text ��� ���  ��� � ����� ��������������� ����������� ������ ���������� -�   ������������� ������������. ���� ��� ���������� ������ �� �  �������� ������ � ��������.!�G /I /Jump /Link f:\work\exper�  t\hlp\login.bmp /Macro /Play /Popup /Just C!�� /P /Just L /�  �1,(Global), 0,<LL1>!�( ������� ����,(Global), 0,<UserInter�  Text � ������������ ������ ����� ����� ������� ������ ���� �  ������ ������ � ������ ������ "OK". ����� ��������� ����� �  �� ����������.!�a/P /Just L /Text ��� �������� ����� ������  ��� ������� ���� ����������. ����� ���� ��� ������ ���������  ���� ����� �������� ������� ������� ����������, �� ������ �    ���� ������ ������  
� �                                 �  /Play /popup /Just L /Text ��������� ������ ���������� �����  � ��� ���, ���� ��� �������� ���������� ������. ���� ������_  � �������� ���������� �������, �� ��� ��������� ������ ����  ��� � ������� P�     �  �� 	`4  �-�   !�* /T N /Just�  cro /Play /Popup /Just C!��/P /Just L /Text � �������������  ������.!�H /I /Jump /Link f:\work\expert\hlp\acc_ch.bmp /Ma�  ���. ���������� ���������� ������ ��� ��������� ������ ����  face>!�" ������ ������,(Global), 0,<(None)>!�! ���_�������,�  �   �&�� 
: # * ?     � Topic@  �    �    �  �    �  ��1N     �  �� 8d     � Topic2�� Gt     � �   �� 	W�   . -�   !�$ /T N /Just M /Text �����������������      
m }                                                     B /Just L /Text ���� ������!� /B /Just L /Text ���� �������  �������:!�* /B /Just L /Text ������������� ���� ������!� /�  ��� ���������� ��������.!�' /S /Just L /Text ��������� �� ��  ����� �� ��������� �������. ���������� ������� � ����� �����  t  x4�� 
� * 1 J     � Topic@Protect  �    �    	  � 2998   �  ��8Y     �  �� C�   *  �% ������ ����    � 2997   �  ��6W     �  �� A~     � ��������� ����   �� ������ ������������� ������� ����� ������� �������� � �    mp /Macro /Play /Popup /Just L  
� �                     �  � ������������!�G /I /Jump /Link f:\work\expert\hlp\acess.b    ���  
� �                                                �  Adm_Users /Link /Macro /Play /popup /Just L /Text ����������  acro /Play /popup /Just L /Text ����������!�K /K /Jump Dlg_�  opup /Just L /Text ������!�H /K /Jump Dlg_Adm_Ergo /Link /M�  � �����������������.!�1 /S /Just L /Text ������ ����� ������  ������� ������� ������� ������ ����� ������ ����� ����� ����  � �� ������ ���������� ��������������.!�` /P /Just L /Text �  ��. ������� ���������� �������� ���������� ���������� ������  ��. �� ����� ���������� ��� ����� ������������� ������ �����  ��� ������. ������ ������������� � ������ ���� ������������  ��� ����� ������������. � ����� ������ ��������� ������ ����  ��������, ������� ����������� ����� ��� ����� ���� � �������  �������� �������. �� ������ ��������, �� ����������� �������  f  O�� 
� . 5 N     � Topic@Dlg_Adm_Acc  �   �  �� ����������. ���� ��� ��������� ����� ���������� ����� ���  ����, �� ������� ���� ���������� ������ ���������� ��������  ��.!�� /B /Just L /Text �������������� ����� ��� ������ - ��  ����� � ��������� �������� ���� ����� ���������������� ����    ������� � ����� ������������ �������.  
� �                 �������� XOR � DES.  
� �                                �  �� ����) ��������������.������� ��������� ���������� ��� ���   ������������� ���������, � ������ (���� ������ �������� ��  �� ������, �� ��� �������� ������� �� ������ "OK" ��� ������  ������ � ������ ������ �� ��� ����������. ���� ��������� ���  ���� � �����, ������ �������� � ����� ���������� ��������� �  ���� �������������� ��������� ������������� ����� ������� ��  N /Just M /Text ������!��/P /Just L /Text ��� �������� ����  �����������.�������� V�     �  �� 	f]  �-�   !� /T �   �  	  � 2996   �  ��<]     �  �� G�     � ������b�  �������� ������, ��������� �������� ���� ���������� � ������  �������� ������������.!�5 /B /Just L /Text ����������� �����   /Text ���������� ������ ������������.!�' /B /Just L /Text �  ����).!�# /P /Just L /Text �������� ��������:!�0 /B /Just L�   ��������� ������� ������������ � ����������� (����� ��� ���  ������� �������������� ������������� ������ ������������� ��  ,  ,��� 
� 0 7 P     � Topic@Dlg_Adm_Users  �  �    �  	  � 2994   �  ��>_     �  �� I�   #  � �����  �������������.�������������� X�     �  �� 	h#  {-�  �   !� /T N /Just M /Text ������������!�� /P /Just L /Text ���  �  Q��� 
� / 6 O     � Topic@Dlg_Adm_Ergo  �  �    �  	  � 2995   �  ��=^     �  �� H�   !  � ������  ������������.������������ W�     �  �� 	g�  -�   !��   /T N /Just M /Text ����������!�T /P /Just L /Text ��������  �� �������������� ����������� ���������� ����� ������ - ����  :!�� /B /Just L /Text ���������� �������� ��� ������ - ����    ������ ������������.  
� �                               �  ��������� ��������� ����� ������� ��������� � �������� � ���  ����� ����� ������.!�1 /S /Just L /Text ������ ����� �������   ������������!�F /I /Jump /Link f:\work\expert\hlp\help.bmp�   /Macro /Play /Popup /Just L!�r/P /Just L /Text ����� �����  ������� ��������� �������� ����� ��� ������ ���������� ����G  �� ������������, ����, ���� ������ ��������� ������, ����� �  �  ��� 
� - 4 M     � Topic@Window_All  �    �  �  	  � 3030   �  ��;\     �  �� F�   ,  �' ��������  ��� MDI ������ ���������� �������� U�     �  �� 	e�  �  -�   !�< /T N /Just M /Text ���������� MDI - ������ ������  ����� ������!�� /P /Just L /Text ����� ���� "���� ����������  � ������" �������� ������� ���������� ��������� MDI-������.3   ��������� ������������� ����� ���� � ������ ������������ �8  V  ��� 
� . 5 N     � Topic@Admin_Admin  �   #    !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !��  ����� ������������� ������������ �������� F1 ��� ������� ���  ����� ����. ���� � �� �������������� ������ � �� ��� �����:  ��, �� ��������� ��������������� ������ � ������� ���������    �� ������ ���������� ������ ������������.  
� �          �  ust L!�[ /P /Just L /Text ��������� ������ �������� ����� ��  p /Link f:\work\expert\hlp\about.bmp /Macro /Play /Popup /J�  =  }��� 
� ( / H     � Topic@Login  �    �  	
  �  �Q�� 
� 2 9 R     � Topic@Admin_ChangeLvl  �       
� �                                                    �  �  �U�� 
� * 1 J     � Topic@HelpHlp  �    �  �  	  � 3040   �  ��8Y     �  �� Cw     � ������� ���  ������ R�     �  �� 	b�  /-�   !�! /T N /Just M /Tex�  t ������� ������!�a/P /Just L /Text ����� ���� "������" ���  ������ ������ ��� �������, �� ����� ������������ ������ �� �  ����������� ������� � ��������� ���������� ������� ������ ��  ���� ������� �������� ������ ��������������� � ������. ��� �  ������ �������� ���� ���������� �������. ������������� ����  �. ������ ��������� ��� �������� ����� �� � � ������ �������  ����� ����� ���� ������� �������, ��� ��������� ��� � �����  st M /Text ����� ����� ��!��/P /Just L /Text ���������� ���  ���� ����� ���� [�     �  �� 	k0  �-�   !�! /T N /Ju�      �  	  � 2993   �  ��Ab     �  �� L�     � ��  9  �"�� 
� 3 : S     � Topic@Dlg_FolderSelect  �      
� �                                                   �  ink f:\work\expert\hlp\exit.bmp /Macro /Play /Popup /Just L�  st L /Text ������ ����� ������ ������������.!�F /I /Jump /L�  � ���� ������ ������� ���������� ������� ������.!�2 /S /Ju�  ��� �������� ���� ����� ��������� ����������� �� ��������� �  �  ̆�� 
� - 4 M     � Topic@File_Close  �    �  �  	  � 3003   �  ��;\     �  �� F~     � ���� ��   ��: ��������� U�     �  �� 	e~  �-�   !�- /T N /Just�   M /Text ������� ���������� �������!�*/P /Just L /Text ���b  ����� �� � ������ �������. � ��������� ������ ����� �� ����  L /Text ��������� ������ �������� ���������� �������.!� /BL    /Just L /Text ����� ������� ����� �� � ������� ���������� �  (Global), 0,<FuncToc>!�1 ������������ ������� ����������,(G    ��� ���������.  
� �                                        ����������� "������" � "������" ������ ����� ��������� ���  � �� �������� ����� ��������� �� ��������� �� ������� ����.  ro /Play /Popup /Just L!�� /P /Just L /Text � ������� �����  �� ������.!�D /I /Jump /Link f:\work\expert\hlp\up.bmp /Mac	  �� �������� ����� � ������������ ����� ����� ����� ��������
  ��� � ������ ���� ��������������� ������� �� ������ �������  L /Text ������ ���� ��������� � ������ �����. ����� ��� ���  ���.!�& /S /Just L /Text ������� ������ �����.!�� /P /Just   �� ����������� ������������� � �������� ���������������� ��  �� ��� ������� ������� ����� ����, ������� ����� �������� �  ���� �� ���������� � ����� ������� ������ � �������� ������  ��" � ������� ���� ������� ������� ������� ��.!�> /B /Just     	  � 3005   �  ��:[     �  �� E�   !  � ��������  � ���������� ��������� T�     �  �� 	ds  �-�   !�/ /  T N /Just M /Text ��������� ���������� �������!�/P /Just   L /Text ���������� ���������� �������. ��������� ������ � �=  ���������� ��. ���� �������� ���� � ������ ������ ���������    k\expert\hlp\new.bmp /Macro /Play /Popup /Just L  
� �     t ������ ����� ������ ������������!�E /I /Jump /Link f:\wor     ���� 
� - 4 M     � Topic@File_NewES  �      �  	  � 3001   �  ��;\     �  �� F�     � �������   ���������� ��������� U�     �  �� 	e  v-�  	 !�3 /T   N /Just M /Text ������� ����� ���������� �������!�� /P /Ju  st L /Text ���������� �������� ����� ���������� �������. ��  ���� �� ����� ���� ������� ������� � ������� ������ �������   ��� � ��������� �����. !�) /S /Just L /Text ����� ��������   ����� ��:!�[ /B /Just L /Text ���������� ������ "����� ���b  |  	��� 
� , 3 L     � Topic@File_Save  �    �{    �  	  � 2999   �  ��>_     �  �� I�     � ����^  �  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�      Just L /Text ����������� �������  
� �                   $  �����������!�L /K /Jump EventSh /Link /Macro /Play /popup /%  .!�A /K /Jump Calc /Link /Macro /Play /popup /Just L /Text &   �������� ������ ������ ������������ � ������������ �������    mf /Macro /Play /Popup /Just L  
u �                     *  n  W��� 
� , 3 L     � Topic@File_Open  �    �+    	  � 3002   �  ��:[     �  �� E�     � ������� ,  ���������� ��������� T�     �  �� 	de  �-�   !�- /T -  N /Just M /Text ������� ���������� �������!�
/P /Just L /T.  ext � ���� ������� ��������� ������� ��� ����� - ����������3   � ��. ��� �������� ������������ �������� ������ ���������� 0  �  ~G�� 
� . 5 N     � Topic@File_Recent  �   *   �  	  � 3006   �  ��<]     �  �� G�   #  � ������"  �  �v�� 
� 0 7 P     � Topic@UserInterface  �  3  ����������� � ����������� ����� C++. � ��� ����� ������� ��4  ��� ����������� ����������. ��������� �������������� ������5  �������� ������ ������������ ��� ���������� ���������.!�( /6  S /Just L /Text ������� ��� ����������:!�l/P /Just L /Text7   -(100.25 - Sqrt( 0.0625 ) + min( 10, min( 20, min( 8, min(8   cos(0), min( 6, min( 5, min( 4,9)))))))) + 101�������: 0 [9  Double]����( 0.5 >= 25/5 ||  !(0.5 >= 25/5) && !1 ) || Cos(:  0) == 1�������: True [Boolean]����Scas( "ABC" + "XX" + "CC";   + "12" + "M",  "CC" )�������: True [Boolean]����integer(Sc<  as( "ABC" + "XX" + "CC" + "12" + 'M',  "M" ) ) + integer(Cm=  pi( "abc", "AbC"))�������: 2 [Integer]����string( min( sin(>  0), max(cos(1), tan(3.14))) ) + "   " + string( max( sqrt(1?  .0/3), sqrt(3.0/1)) )�������: 0,000000   1,732051 [String]�@  ���(bbs=1.0) + pow( 2,  9/3*sqrt(9)/sqrt(sqrt(81)) )�������    : 9 [Double]��  
z �                                     b2  ����� LL(1) ����������� � ��������� ��������� ��������� � �F  � ���������!� /S /Just L /Text ���������!��/P /Just L /Te    ��� ��������  
z �                                       C  usLine /Link /Macro /Play /popup /Just L /Text ������������B  p Grammar /Link /Macro /Play /popup /Just L /Text ���������^  xt ��������� � ������� ���������� � ���������:�����������_�    �� ������ ���������.   
� �                              G  ����������� ������ ������� � ��������� ���� � ������� �����H   /Text ����������� �������!�m /P /Just L /Text ��������� ��I  � ��������� R�     �  �� 	b8  � -�   !�& /T N /Just MJ  	  � 2991   �  ��8Y     �  �� C|     � ����������K  A  ���� 
 * 1 J     � Topic@EventSh  �    �  N  t  T��� 
 ' . G     �
 Topic@Calc  �    �  	 O   � 2992   �  ��5V     �  �� @q     � ������������P  � O�     �  �� 	_k  �-�   !� /T N /Just M /Text ����A  �������!�/P /Just L /Text ������� �� �������������� �����`  � 2990   �  ��4U     �  �� ?�   %  �  ���������, ���a  _��������� = ��.������������� = <��1|�������1, [������], [�R  - "������1" + "������2"������� ��������� ���������  �������S  ��- ���_����������1 <= ���_����������2��- !���_���������鑒T  + 55��- ���_����������1��- 55��- -55��- ���_���������� - 10U    ��- ���_����������1 * ���_����������2��- ���_����������1 V  ���� �������� ��� �������) � '!'(������ ������).��������:  W  >=,==,!=}. ��� ��� ��������. ���������� �������� '-'(����� X  �� �� � �����.���������� = {+,-,*,/,%}; {||,&&,!}; {<,>,=<,Y  � ������ ������� � ��� ������ ���������� � ����� ��� {_,@} Z  ��������� = {A..Z, a..z, 0..9, _, @}. ��� ��� ����� �� ����[  �����(5.5); ����������(true/false); ����-��("���"). �����_�\  ��������]>, ���:���ONST = ������('A'); �����(55); ���������]  �������� = <CONST|���_����������1, [CONST|���_����������2, E  N /Just M /Text ���������, �������������� ������!�M /K /Jum_  ����������� �������� N�     �  �� 	^W   �-�   !�3 /T bp  �2|�������2, [������], ��������1, ��3|�������3, ��������2, q  ��� -,*,% � / �� ����������� ��� ��������� ����������). ���b   ����� ��������� ����������� ����� ��� ������� � ��� (�����c   double � ��������� ����� ����� ���� ��� ). ������ ��������d  ��� ���������� (5.0 + 2 - ����� ��������� ����� ��������� �e  ��� ���������� ����� ����������� � ��-��� ������� ���� �� �f  (ABC))) ).��������� ���� �� �����������. ��� �������� �����g  �����" || !ABC || Min(C1, C2) > 2��- Cos( Sin(X*C - Tan(Cosh  (C * C) || (B2 > 0)��- A1 + Cos(C * C) || B2��- Start@ == "i  �������2 + ���_����������3 < 2��- A + (C - D)/2��- A1 + Cosj   ���_����������. ��������:    ��- ���_����������1 * ���_���k  ouble,string}-���������� ����� ������ ���.�������_������� =l  qrt,floor,ceil,exp}-������ ����-�����. {bool,char,integer,dm  ��� ����������. {sin,cos,tan,atan,asin,acos,log,log10,exp,sn  ���������1, [���������2]). {min,max,pow,fmod,cmpi,scas} - �o  .., ��N|�������N, ��������N]>, ���:��������� = ���_�������(b�  ���� ���� ����� ����������� �� ����. ��������� ������� (min�  ����������� ������.��-����� - �����. ������� ���������� - �r  ������ ���� �� ����������� � �������� ������ � ���������� �s   �� ���������� �������� ������� ������. ����� ���������� ��t  �������� ��� ���������� ����������). � ���� ������ ��������u  ������ ����������, �������� � ������� (������� ��������� - v  ���� ������� - ����������� ��� ������������ ������������� �w  � ������������ 0-1)!��/P /Just L /Text -����� - �����. ���x  ����.!�E /S /Just L /Text ������������ ������� (�����������y  ��� �������� ����������. ����� ������ �� ����������� ������z   � ���������� ����������� � ����� ����� ������ ���� �������{   ����� ��� A + B, �� ����� ������������� � ���� bool(A+B)).|  � ����������� ���������� ���� � bool (�������� ���� �������}  �� ���� (sin - ������ double).����� ��������� ������� �����~  ���������. ������ ������� ���������� ��������� ������������  , max) ���������� ��������� �������� ������� ���� �� ���� �  ���������� ��������� ��� ������ ����� ������� 100% ������. �  ��� ������ ������� �������� � ������ ���������� ������������  (B|A)= P(B)*P(A|B) - �������� ���������������� ������ ���� �  B)- P(A)*P(B) - ��� ��������� ������鑒(4)  P(A*B) = P(A)*P�  �� ������������� ����������� ������鑒(3)  P(A+B) = P(A)+P(�  ������鑒(2)  P(A*B) = P(A)*P(B) - ����������� �������������  1)  P(A+B) = P(A)+P(B) - ����������� ������ �� ����������� �  ��� ������.��� ������ ������ ���������� �������� ������:��(�  �� ������ � ��� �������� ��� ��� ��� ����� ������ �� �������  �������� ��������� �� ���� ��������� ��������, ������� �����  ���, �� ���� ����� max. � ����� ������� ������������ �������  ����� ���������� ��������� �. ���� ��� ��������� ��������� �  ��� ����������� ��� ������� ���������, ��� N ������� �������  �������: ����� = �����*min( �����1, ..., �����N) - ��� �����  ��������� �������� � ���������� ���������-��� �������. �����  ��-����� - �����. ������� ������ - ����������� ���������� �    ������� ������ ������ ��-��� ����������� �� ������� (3). (�  1_2; �������2;..; �������N �� ����������1, ����������1_2:���  ����� ���������!��/P /Just L /Text ����  �������1, ��������  ��������� 2,.., ��������� N )* ����.!�" /S /Just L /Text ���  ������ �������� ��� "�", ����� �������� = min(��������� 1, �   ����������1, ����������2,.., ����������N :����   - ����� ��  ������1* ����.��������  �������1, �������2,.., �������N  ���  ��1, ����������2,.., ����������N  :�����   - �������� = ����  � 2,.., ��������� N )* �����.��������  �������1 �� ���������  ������ ��� "�", ��-��� �������� = min(��������� 1, ���������  �2,.., �������N  �� ����������1  : ����� - ����� ������� ���  � - �������� = ���������1* �����.��������  �������1, �������  .!�2/P /Just L /Text ����  �������1 �� ����������1  : �����  ����������� �� (3))��!�# /S /Just L /Text ������� ����������  ���������� ��-��������, �� ����� �����. ������� ���������� �  �� ���� ���� ���� ����� �������� ������������� ��� �������肰  ���1; �����-�����2:�����2;..; ����������N:�����N   - ����� �  �� ���������.!�% /S /Just L /Text ���������� ���������!��/�  �� ���������� �������� � � ������ ������������ ������ ������  ��� ��������� � ������� � ����������, ������������� � ������  �����. ������ ��������, ��������� ������������ ������ ������   �����-����).������ ���������� ����������� �� ������� ������  � ��� ����� ���������� ��� � ����� ���� (����� ���������� ��  ����. ��� ��������-����� ������� ��������� ������� ���������  ��� � �������� ����� ���� � �� - ������ ��� ������� ��������   ���������� ����� �������, �������-���, �� ��������� �������  ��������:  ����� ��������� ����� ����� ��������. �����������  �- ���� A>2, CS=="�����" �� M = Cos(Min(A-B, C)) :0.9�������  �>������ = ��������� ���������������������� ���������:    ��  ��� = ��������ő����������� = <���_����������,  =, ���������  � ����������� �� ��������� "���" (����� � �������).���������  ��������� ����������� �� ������� ��������� �������������-����  P /Just L /Text � �������� � ����������� ��������� ���������  ������ {True, False};��- ����� ��������� {10};��- ����������  �� ������� - �������. ��������� ��������:��- ���������� ����  �������� ������� ������� ������������ �������� �� ����������  /Popup /Just C!�|/P /Just L /Text ����������� ���������� ��  �F /I /Jump /Link f:\work\expert\hlp\synt.wmf /Macro /Play �  �����  � ������ ���������� ������� �������� ��� ���������.!�  �� �����.������ ������� ��������� - ���������� ������ ��� ��  ������� �������� ��������� � �������������� ������ ���������  �� ������ � ���������� ������ ������ ��� ���������;��- ����   �� ��� ������:��- ���������� LL(1) ����������;��- ��������   "=". ������ ����������� ���. ����������� ��������� ��������  �� ������ ��������� �� ����� � �� ����� ������ �������������  ���������� "=". �� ���������� �������-������ ���������� - ��  ���� ������������� ����������� - ��� �� ������ ��������� ���  ���� ��������� ��������������� ���������� ����� "C". �� ����  ����� ��������� � ������������� ������ {7.25};��- ����������  ���� �����. ������� ����������� ������ ������, ������� �����  ���������� �� ������� ������ ����������� ����������� �������  ������� ���������� ���������� ���� ������. �� ��������� ����  ��-�� ������ �������� ���������� �� ���� �������. ����������  ���� - �������������� ���������, � ������ - ��������� �� ���  �� ��������� ���� <���_�������, ������>. ������ ���������� �  �� - ��� ������� ������������ ��������, � ������� ����������  � ������� � ������ ���-����������� ������� - �������. ������  ������� � ���, ����� ������������� ����������� ������������  ��- ������� ������ {(, )};��- ������� {,}.����� ������ �����  ����� �������� {*, /, %, +, -};��- �������� ���������� {=};�  ;��- ������������� {���_����������, Sin, Cos};��- ����������  };��- ���������� �������� {||, &&, ==, !=, >=, <=, >, <, !}�  ��������� ��������� {'C'};��- ��������� ��������� {"������"�  ����� ��������� � ��������� ������ {0.25E+15, 0.8E-5};��- �b�  �������� ������-�������� ��������� ���������. ���� ������ ��  �����.!�p/P /Just L /Text ��� ���������� ��������� ��������  � ��� ��������� �� ��������� �� �������. � ������ ����������  ���� ��� ��� �������� ���������� ������ ����� �� ��������� �  ������� � ����������� ������� ������ ������� ����. ��� �����  ��� ��� �������� ����� ������� ���� ����� ��������� ������     ro /Play /Popup /Just L  
� �                            �  � ������:!�E /I /Jump /Link f:\work\expert\hlp\ll1.wmf /Mac�  Sin(1) + min(2, Var3)*2) + 10.5) / pow(2, 3) �������� ������   /Just L /Text ��� ���������� ��������� (Var1 + 25/Var2 - (�   ����.!�+ /S /Just L /Text ������ ������ �����������:!�� /P  ��,(Global), 0,<Exp_Pane>!� ���������,(Global), 0,<LL1>!�+�  lobal), 0,<LL1>!� �������,(Global), 0,<Explorer>!� �������   ����� ��������� ��������, ���� ���������� ����� ��� �������  ����� ������ ������� ���� ������������ ���������, � ��������  ����������� �� ��������, ������� ���� ���������. ������ ��-b�  �� ��� ������, ��� ��������, ��� ������, ������ ��������/���  ��� �������� ������� ����. �� ����� ���������� � ������� ���  /Just L /Text ������ ������� ��.!�b /P /Just L /Text �������  k\expert\hlp\exp_imp.bmp /Macro /Play /Popup /Just L!�# /S �  �������� ��������������� ��������.!�I /I /Jump /Link f:\wor�  .!�� /P /Just L /Text � ����������� �� ��������� ������ ����  opup /Just L!�, /S /Just L /Text �������� ������ ������� ���  /I /Jump /Link f:\work\expert\hlp\e_new.bmp /Macro /Play /P�  �4 /T N /Just M /Text ������ ������������ ���������� ��!�G     ext ������� ����  
� �                                   �  �� �������� ��� ������������� ����. ����� �������� ����� ���  �� ������ ������������� ���� ������ ��� ���� ������ ��� ���  �  ���� 
� , 3 L     � Topic@Work_Pane  �    �|   � 3986   �  ��5V     �  �� @�      � ������ �������  ust C!�� /P /Just L /Text ����� ��������� �� ����������� ���  � ��������� ���������� ������: ��������� �����, �����������   ����� ������ ��.!�I /I /Jump /Link f:\work\expert\hlp\exp_r�  }
  ��� 
� + 2 K     � Topic@Exp_Pane  �    � �   	  � 2988   �  ��9Z     �  �� D�   &  �! ������ ���  ���������� ���������� ���� S�     �  �� 	ct
  �	-�   !  �� ������� (�������) � �������� �� � ������/������ ������� �  ext ������ ��������� �������� ��.!�] /P /Just L /Text ������  lp\exp_uns.bmp /Macro /Play /Popup /Just L!�. /S /Just L /T�  ��� ������������� �����.!�I /I /Jump /Link f:\work\expert\h�  ��������, ���� �������� ����, �� ��� �� ����� ������ ������  ��������� �� �������� ��������� �������� �������� �������. �  L /Text �������������� ������� ��.!�� /P /Just L /Text � ���  ert\hlp\exp_ed.bmp /Macro /Play /Popup /Just L!�+ /S /Just �  ��� ������ �� ����������� ��.!�H /I /Jump /Link f:\work\exp�  ��. ����������� ������� ��������: � ������ ������� ���� ����  ���� ������� ��.!� /P /Just L /Text ��������� ������� �����  em.bmp /Macro /Play /Popup /Just L!�% /S /Just L /Text ����b�  Link f:\work\expert\hlp\exp_tree.bmp /Macro /Play /Popup /J  ��������� ���� �������� ��.!�? /P /Just L /Text ������� ���  bmp /Macro /Play /Popup /Just L!�3 /S /Just L /Text ������   ����� �����.!�J /I /Jump /Link f:\work\expert\hlp\exp_uall.0   ������������� �������,(Global), 0,<Protect>!�# �����������  <  b#�� 
� + 2 K     � Topic@Explorer  �    �    	  � 2989   �  ��9Z     �  �� Dv     � ���������	   ���� S�     �  �� 	c3  �-�   !�. /T N /Just M /Text
   ��������� ���������� ������!��/P /Just L /Text ����������   ��������� ���������� ������� � ��������� ������������� �   ��������� ���������� � ��������� ��� ���� ��������������� �  �������. � ���� ���������� ��� ������ � ���� ������. ������   �������� ������������� ���� ������ �������, � ���� �������  , �������� ������ �������� � ������. ���������� ��� ������   �������� ������������� ���� � ������. ������� ����������� �  ������������� ��������� � ������������� ����.!�J /I /Jump /�   ���� (�������) �� ���� �������� ��.!�I /I /Jump /Link f:\wo!  �� ���������� ������������� ���� ������. ����������� ������  !�� /P /Just L /Text �������� ������ ������������/������� �  acro /Play /Popup /Just L!� /S /Just L /Text ������������.  � ������.!�G /I /Jump /Link f:\work\expert\hlp\exp_q.bmp /M  ust L /Text ����������� ���������� ���� � ������������� ���  L /Text ���������� ���������� ������������� �����.!�I /P /J  t\hlp\exp_comp.bmp /Macro /Play /Popup /Just L!�; /S /Just   �������� ������� � �������.!�J /I /Jump /Link f:\work\exper  �������� ������ ��������������. ��������� ������� ������ ��  /Text �������� ������ ��������� ���� ������� � ������� ��.   t L!�% /S /Just L /Text ������ � ������� ��.!�� /P /Just L   ink f:\work\expert\hlp\exp_sec.bmp /Macro /Play /Popup /Jus  � ������ ��������� ���������� ���������� ��.!�I /I /Jump /L   /Just L /Text ��������� �����.!�D /P /Just L /Text �������  rk\expert\hlp\exp_opt.bmp /Macro /Play /Popup /Just L!�! /Sb    � ���� �������� � ������.  
� �                          1   �������� �������� ��� ������ ����, �� ����������� ��������"  �� ��������� ����� C++. ���������� ����� ����������. ���� �#  /P /Just L /Text ��������� ��������� ������������� ��������$  ����� ������ ���������. �� - �������������� ����� 0..1.!�&%  �� ������������. � ��������� ����� ���� � �� �� ����� - ���&  �� ����������� - ������ ��������� ���� � ������ ���� ������'   ������ ��������� ������������. �� "���������2" �����������(  ��������2 :��>���� "���������1" ������������� ����������� -)   ������ ���������!�I/P /Just L /Text <���� ���������1 �� �*  � �������������� ��� ������ � ��������.!�! /S /Just L /Text+   ������� ��������������� �����������. ������������ ����� ��,  ��������� � ����� ������. ��������� ������������ �� ����� �9   L /Text ��������!�0 /P /Just L /Text ������� ������� �����.  ert\hlp\exp_uns.bmp /Macro /Play /Popup /Just L!� /S /Justr  ,(Global), 0,<Work_Pane>!�( ���������� �������,(Global), 0,�@  �� � ����� �������� ���� � ��������� ����� ����� ����. ����A  Text �������� ��������� ����� ���������� ���������� ���� ��2  /Popup /Just L!� /S /Just L /Text ��������!�L /P /Just L /3  I /Jump /Link f:\work\expert\hlp\pro_uncm.bmp /Macro /Play 4  �3 /P /Just L /Text ��������� ��������� � ���� ������.!�J /5   /Macro /Play /Popup /Just L!� /S /Just L /Text ���������!/  ������ �� ������������� ����.!�I /I /Jump /Link f:\work\exp7  ext ������ ���� ������!�> /P /Just L /Text ��������� ������6  � �� ����.!�I /I /Jump /Link f:\work\expert\hlp\pro_cmm.bmp]  ������, ������������ �������>!�h /P /Just L /Text ���������:   /Just L /Text ������ �������!�7 /P /Just L /Text <���_����;  ��� = �������� :��>���������� ������ ���� ����������.!� /S<  /Just L /Text ������ �����!�R /P /Just L /Text <���_�������=   �������������� �������, ������������� Visual Expert!� /S >  �l /K /Jump FuncToc /Link /Macro /Play /popup /Just L /Text?  ���� ��� �������� integer � double ��������� ����� double.!�P  ����.!�J /I /Jump /Link f:\work\expert\hlp\exp_comp.bmp /MaC  ���������� ��������� ������������� ����� S�     �  �� 	D  c=  �-�   !�B /T N /Just M /Text ������ ������������ ���E  ������ ������������� ���!�I /I /Jump /Link f:\work\expert\h8  lp\pro_rdc.bmp /Macro /Play /Popup /Just L!�# /S /Just L /T     ������.  
� �                                           F  xt �����!�7 /P /Just L /Text ������� � ��������� ����������G  \pro_exit.bmp /Macro /Play /Popup /Just L!� /S /Just L /TeH  ����� ����� ���������.!�J /I /Jump /Link f:\work\expert\hlpI  /Just L /Text �����!�: /P /Just L /Text ������� ������ ����J  k\expert\hlp\exp_opt.bmp /Macro /Play /Popup /Just L!� /S K  �������� ���� ����� � ���� ������.!�I /I /Jump /Link f:\worL  pup /Just L!� /S /Just L /Text �����!�4 /P /Just L /Text �M  /Jump /Link f:\work\expert\hlp\pro_sch.bmp /Macro /Play /PoN  �1 /P /Just L /Text ������������ ������ ���� ������.!�I /I O  cro /Play /Popup /Just L!� /S /Just L /Text �������������!�B   	  � 3987   �  ��9Z     �  �� D�   4  �/ ������ ��a  ������ �������� ���������� ������� ���������� ����:!�9 /B /R  t ����������� ���� ����������!�M /P /Just L /Text ��� �����S  /Play /popup /Just L /Text ������ ������!�, /S /Just L /TexT  ���� ������� ����������.!�G /K /Jump Tree_Res /Link /Macro U  ������ �������� ������ ��������������� �� �������� ��������V  ��������� ����� ���� ���������� �� �������� � ����� ��������  � ����������,(Global), 0,<Protect>!� ������,(Global), 0,<PZ  � ���������. �� ���� ��������� ����������� ������ ������ ��[  ���� ������� ����� ������������. ������ ������ ��������� ��W  � �������� ������ � ��������� �������� ��������� �������.���  �� ����� ���������.!�W /K /Jump Pro_pane /Link /Macro /Play\   ����� ��������� ������ � �������� �������� � �������������  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�   �� Visual Expert!�Q /L /Jump HotKeys /Link /Macro /Play /poQ  F  L�� 
F + 2 K     � Topic@Pro_pane  �    � 6p  Just L /Text ������������������ ���������� (�������).!�B /Bq  � ������������ � ��������.!�U /K /Jump Work_Pane /Link /Macb  ������.!�J /P /Just L /Text � ��������� ���� ������� ������c  st L /Text � ��������� ������.!�  /B /Just L /Text ����� ��d   ������ ����� �� ������������ - ������ ���������.!�$ /B /Jue  ����� � ��� �������:!�S /B /Just L /Text ��� ������� - ���f   ������ ������ ������ ������!�0 /P /Just L /Text �������� �g  /Text ������� - �������������� �������.!�, /S /Just L /Texth  ���� ������� - ��������� ������������������.!�2 /B /Just L i  ������ ��������� ������� ���������.!�@ /B /Just L /Text ���j   /Just L /Text ���� ���������!�= /B /Just L /Text ������� �k  ��� � ������� ������ ����������� �������� ����������.!� /Sl   /Just L /Text ��������� �� ������� ������ ����� �������� �m  �2 /B /Just L /Text �� ������������������ ����������.!�r /Pn  ���).!�1 /B /Just L /Text ��������� ���������� (�������).!o   /Just L /Text ���������� �� ����� ��� ����������� ���� (�肀  ro /Play /popup /Just L /Text ������ ������������ ������  u  <Protect>!�= �������������� ���������� LL(1) �����������,(Gt  ������� ��� ��������� ����������. ������� � ������ � ������  ����� ������ ��������� � ������� ����������. ����� ���� ���X  lobal), 0,<LL1>!� ������,(Global), 0,<CreNewObj>!�' ������  ������ S�     �  �� 	c�  �-�   !�  /T N /Just M /Texv   	  � 3984   �  ��9Z     �  �� Dw     � ������ ��w  �  �?�� 
r + 2 K     � Topic@Tree_Res  �    � Y  ����� � ��������� ������������ ������� ������ (���� �����) y   ��������� ��������� ������ ������ ��� ������������� ���� �z  ust M /Text ������ ������������/�������!��/P /Just L /Text{  ������/��������� O�     �  �� 	_Y  �-�   !�. /T N /J�  !�- /B /Just L /Text ������ ������� - ����������.!�0 /B /Ju}  ���������� ����.!�' /S /Just L /Text � ������ ������������:~  �������� - ����� �������� � ��������������� �� �������� ��     
� �                                                      b    ��� ������� ������� � �� � �������� �����.  
� �         �  ext �����/����������!�2 /P /Just L /Text �������� ������ ���  ������� ������.!�J /I /Jump /Link f:\work\expert\hlp\pro_ex�  it.bmp /Macro /Play /Popup /Just L!� /S /Just L /Text �����  �!�( /P /Just L /Text ������� � ��������� ��.!�H /I /Jump /�  Link f:\work\expert\hlp\w_stop.bmp /Macro /Play /Popup /Jus�  t L!�# /S /Just L /Text ������� (Shift+F5)!�" /P /Just L /T�  ext ���������� �����.!�G /I /Jump /Link f:\work\expert\hlp\�  w_prt.bmp /Macro /Play /Popup /Just L!� /S /Just L /Text �s  .bmp /Macro /Play /Popup /Just C!�� /P /Just L /Text �������  t ������ ������!�H /I /Jump /Link f:\work\expert\hlp\tree_w�  �����!�H /P /Just L /Text �������� ���������� - ������� �� �  ������� ������ ������.!�G /K /Jump Tree_Res /Link /Macro /P�  lay /popup /Just L /Text ������ ������!�G /I /Jump /Link f:�  \work\expert\hlp\w_ask.bmp /Macro /Play /Popup /Just L!� /�  S /Just L /Text ������!�K /P /Just L /Text �������� ������ ��  lp\exp_opt.bmp /Macro /Play /Popup /Just L!�! /S /Just L /T�  st L /Text ��������������� ������ - �����.!�$ /B /Just L /T�    	  � 3985   �  ��:[     �  �� E�   ,  �' ������ ��  ����������� ������ �������������� T�     �  �� 	d�  (�  -�   !�: /T N /Just M /Text ������ ������������ ������ ����  ���������!�G /I /Jump /Link f:\work\expert\hlp\w_stm.bmp /M�  acro /Play /Popup /Just L!� /S /Just L /Text ������� ������  !�0 /P /Just L /Text �������� ������� ����� �������.!�H /I �  /Jump /Link f:\work\expert\hlp\w_anim.bmp /Macro /Play /Pop�  up /Just L!�& /S /Just L /Text ����� �������� ������!�� /P �  /Just L /Text �������� ����� �������� ������ - ������ ������  � �������� � ����������� ������ � ���������� ���������� �� �  ������ ����.!�H /I /Jump /Link f:\work\expert\hlp\w_step.bm�  p /Macro /Play /Popup /Just L!�! /S /Just L /Text ��� ������  � (F10)!�H /P /Just L /Text ��������� ��� ������ - ����� ���  ������ � ������� ������.!�I /I /Jump /Link f:\work\expert\hb�  ext �������� - �������.!�J /S /Just L /Text � ����������� ��  �� ������ ���� ����� ��� ���� ���������, �� ������ �����. ��  ��� ��������� ��������� ��. ������ ���� ��������� ����� ����  Just L /Text � ������� ����� �������� ����� � ������ �������   /T N /Just M /Text ��������� ����� ������ ��������!�/P /�   ����� ������ ���������� S�     �  �� 	c�  [-�   !�2�   	  � 3983   �  ��9Z     �  �� D�   $  � ����������    ���� 
� + 2 K     � Topic@Work_Opt  �    � �  ���� ����� ������� ������ �������� ������ ������� ������ ���   L /Text �������� � ������ ����. ��� ������ ���� ������ � ��  ���������.!�7 /S /Just L /Text ����� ������� ������������� �  ���� ����:!�O /P /Just L /Text �������� � ������ ����� ����    ����� ������ �� < 0.33.  
� �                            �  �� - ������� 0.67 < �� >= 0.33.!�/ /B /Just L /Text ����-���  ext ������ - ������� �� >= 0.67.!�5 /B /Just L /Text ������  � ������������ ������� ������������ �����:!�. /B /Just L /Tb�  ������ ������ "�����" ����� ��������� ��� ���� ��������� ���  /Text � ����������� �� �������� ������ ����� ��� ������ ����  � ������� �������� ������ � �������� �������� ������� ��. ��  ������� ����� ��������� ��������� �� �������������� ��������  ���� ������������� ��� ������������ �������. ����� ���������   ������ ��� ������� ����� ����� �������. ������� ������ ����  ��� - ���� ����� ������ ����������� � ������� �������� ��.!�  �> /S /Just L /Text ����� ������� ������������� ���� �������   ����:!�Z /P /Just L /Text �������� � ������ ��� ������ ����   ������ � ������ ������ �������� �������.!�+ /S /Just L /Te�  xt ����� ������� ���� ������:!�� /P /Just L /Text �������� �  � ������ ����. ��� ������ ���� ������ � ����� ����� ��������   ������ �������� ������ ������� ������ �����������.!�3 /S /�  Just L /Text ����� ������� ����  �������� ����:!�� /P /Just    � ������ � ������ ������ ��������.  
� �                     ��� ������ - ��������� ��������� ��� �����.  
� �        ��   N /Just M /Text ��� ������� ����� ������ ��!�l/P /Just L �  ������ �������� ���������� � ����� ������� ����. ��-������ �  ���� ������������ ����� � ��������������, �� ����� ���������  � �� ���� ���������� � ��������������� � ��������� ����� ���  Just C!�F /I /Jump /Link f:\work\expert\hlp\tbl4.wmf /Macro�  ump /Link f:\work\expert\hlp\tbl3.wmf /Macro /Play /Popup /�  rk\expert\hlp\tbl2.wmf /Macro /Play /Popup /Just C!�F /I /J�  bl1.wmf /Macro /Play /Popup /Just C!�F /I /Jump /Link f:\wo  A   ��  � ) 	4       � Topic@Topic2	  � 3980   �  b  ��� 
� ' . G     �
 Topic@Work  �    �  	      /Play /Popup /Just C  
� �                              �  ������������� ����. !�F /I /Jump /Link f:\work\expert\hlp\t�  rotect>!� �������,(Global), 0,<FuncToc>!�  !�  !�  !�  !� �  �  O�� 
� , 3 L     � Topic@CreNewObj  �    ��    	  � 3982   �  ��:[     �  �� E�      � ��� �����  ��� ����� ������ ���� T�     �  �� 	d�  T-�  
 !�. /T6�   /Just L /Text ���� ���������� ������� ���� ���������� � ��Q  `   Q��� 
� & - F     �	 Topic@LL1  �    �  	  �   ���������� ��������� ������������ ������ ������ �����������  	  � 3980   �  ��8Y     �  �� C�   8  �3 �����������  ���� �������, ������������� Visual Expert�� R�     �  ��  � 	b�  �-�   !�F /T N /Just M /Text �������������� ������  ��, ������������� Visual Expert!�M /K /Jump Grammar /Link /                                                               �   /popup /Just L /Text ������ ������������ ���������  
� �     !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�        �  q  �3�� 
� . 5 N     � Topic@ProductEdit  �   �   �  	  � 3988   �  ��<]     �  �� G�   &  �! �������  �� ������������� ��� �������� V�     �  �� 	fh  �-�  �   !�4 /T N /Just M /Text �������� ������������� ��� ������!-  �� /P /Just L /Text ������������ �������������� ��������� ��  Macro /Play /popup /Just L /Text ���������� ���������!�/P�    � Topic4                                                 �  '����%right  '!'����%left   '('����/*----------------------�  EQ     GEQ��%left   '+'     '-'��%left   '*'     '/'     '%�    OROR��%left   ANDAND��%left   EQU��%left   NEQ��%left   L�   ANDAND  EQU     NEQ     LEQ     GEQ��%right  '='����%left �         STRING_CONSTANT��%token  IDENTIFIER��%token  OROR   �  AT_CONSTANT  INTEGER_CONSTANT��               BOOL_CONSTANT�  � LL(1) ����������.�� �� �� %token  CHARACTER_CONSTANT  FLO�  ���� ���������. ��� ���������� ������ ����������� ����������  �� ������� ������ ����� �� ������� (Expression), �����������  �	  wE�� 
� * 1 J     � Topic@Grammar  �    �  �  	  � 3979   �  ��8Y     �  �� C}     � �����������   ����������� R�     �  �� 	b�	  	-�   !�' /T N /Just �  M /Text ���������� ���������!�> /K /Jump LL1 /Link /Macro /�  Play /popup /Just L /Text ���������!��/M /Just L /Text ����  A   �  � ) 	4       � Topic@Topic4	  � 3979   �   ----- start symbol ------------------------------*/����%sta  xpression '-' Multiplica-tive_Expression��;����Multiplicati�  ive_Expression '+' Multiplica-tive_Expression��| Additive_E�  ��Additive_Expression��: Multiplicative_Expression��| Addit�  ssion��| Relational_Expression GEQ Additive_Expression��;���  tive_Expression��| Relational_Expression LEQ Additive_Expre�  n '<' Additive_Expression��| Relational_Expression '>' Addi�  l_Expression��: Additive_Expression��| Relational_Expressio�  uality_Expression NEQ Relational_Expression��;����Relationa�  sion��| Equality_Expression EQU Relational_Expression��| Eq�  y_Expression��;����Equality_Expression��: Relational_Expres�  uality_Expression��| Boolean_AND_Expression ANDAND Equal-it�   Boo-lean_AND_Expression��;����Boolean_AND_Expression��: Eq�  ion��: Boolean_AND_Expression��| Boolean_OR_Expression OROR�  �| Unary_Expression '=' Expression��;����Boolean_OR_Express�  rt Expression����%%����Expression��: Boolean_OR_Expression��  ve_Expression��: Unary_Expression��| Multiplicative_Express                                                               D  pup /Just L /Text ������� �������� �������!�T /L /Jump Stat     !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�                �  �  1�� 
� * 1 J     � Topic@FuncToc  �    �      �%%��  
� �                                                T��| FLOAT_CONSTANT��| BOOL_CONSTANT��| STRING_CONSTANT��;�  ion��;����Constant��: INTEGER_CONSTANT��| CHARACTER_CONSTAN  ���Argument_List��: Expression��| Argument_List ',' Express	  ression��: IDENTIFIER��| Constant��| '(' Expression ')'��;�
  ostfix_Expression '(' Argument_List ')'  ��;����Primary_Exp  '!'��;����Postfix_Expression��  : Primary_Expression��  | P  y_operator Unary_Expression��;����Unary_operator��: '-'��|   ession��;����Unary_Expression��: Postfix_Expression��| Unar  nary_Expression��| Multiplicative_Expression '%' Unary_Expr  ion '*' Unary_Expression��| Multiplicative_Expression '/' U